module main

pub fn mgeaprint()
{
	println('Hi this is from mega')
}