module encx

pub fn myprint()
{
	println('Hi, this is from base encode')
}

pub fn extra()
{
	println('Hi, this is from base encode')
}
