module main

fn test_get_totp() {
	key := [u8(0x31), 0x32, 0x33, 0x34, 0x35, 0x36, 0x37, 0x38, 0x39, 0x30, 0x31, 0x32, 0x33, 0x34,
		0x35, 0x36, 0x37, 0x38, 0x39, 0x30]

	data_test := [u64(0x1), 0x23523EC, 0x23523ED, 0x273EF07, 0x3F940AA, 0x27BC86AA]
	result_test := [287082, 081804, 050471, 005924, 279037, 353130]

	for i, item in data_test {
		data :=convert_u64_to_u8(item)
		otp := get_totp(key, data)

		assert otp == result_test[i]
	}
}
